module sobel_g_assertions (
    input  logic                  clk,
    input  logic                  rst,
    input  logic [COLORDEPTH-1:0] vect_in [M_DEPTH-1:0],
    input  logic [COLORDEPTH-1:0] conv_o,
    input  logic                  dv_i,
    input  logic                  hs_i,
    input  logic                  vs_i,
    input  logic                  line_end_o,
    input  logic                  hs_o,
    input  logic                  vs_o,
    input  logic                  dv_o
);


endmodule
