module sobel_top_assertions (
    input  logic        clk,
    input  logic        rst,
    input  logic        h_pol,
    input  logic        v_pol,
    input  logic  [7:0] sw,
    input  logic  [7:0] red_i,
    input  logic  [7:0] green_i,
    input  logic  [7:0] blue_i,
    input  logic        dv_i,
    input  logic        hs_i,
    input  logic        vs_i,
    input  logic  [7:0] red_o,
    input  logic  [7:0] green_o,
    input  logic  [7:0] blue_o,
    input  logic        dv_o,
    input  logic        hs_o,
    input  logic        vs_o,
    input  logic        hs_o,
    input  logic        vs_o,
);

endmodule